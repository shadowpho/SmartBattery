** Profile: "SCHEMATIC1-abc"  [ C:\Users\aaa bbb\Documents\KiCadProj\SmartBattery\pSpice\Design1-PSpiceFiles\SCHEMATIC1\abc.sim ] 

** Creating circuit file "abc.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpiceTIPSpice_Install\17.4.0\PSpice.ini file:
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 30m 1m 
.OPTIONS ADVCONV
.OPTIONS THREADS= 20
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
